.MODEL NMOS NMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 4.1E-9
+XJ      = 1E-7           NCH     = 2.3549E17      VTH0    = 0.3729594
+K1      = 0.5840975      K2      = 1.686187E-3    K3      = 1E-3
+K3B     = 0.0296594      W0      = 1E-7           NLX     = 1.542817E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 1.1680674      DVT1    = 0.4182499      DVT2    = 0.0268331
+U0      = 292.3966054    UA      = -1.219746E-9   UB      = 2.307456E-18
+UC      = 6.953926E-11   VSAT    = 1.704188E5     A0      = 1.8603725
+AGS     = 0.4358979      B0      = 1.843628E-7    B1      = 5E-6
+KETA    = -0.011523      A1      = 8.967934E-4    A2      = 0.3
+RDSW    = 105.3073514    PRWG    = 0.489299       PRWB    = -0.2
+WR      = 1              WINT    = 0              LINT    = 1.963253E-8
+         DWG     = -5.54717E-9
+DWB     = -1.072339E-8   VOFF    = -0.0948017     NFACTOR = 2.1860065
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 1.925032E-3    ETAB    = 6.028975E-5
+DSUB    = 0.0193048      PCLM    = 1.9022344      PDIBLC1 = 0.2550871
+PDIBLC2 = 1.417207E-3    PDIBLCB = -0.1           DROUT   = 0.8645309
+PSCBE1  = 3.419362E10    PSCBE2  = 2.777738E-8    PVAG    = 9.459578E-3
+DELTA   = 0.01           RSH     = 7              MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 8.58E-10       CGSO    = 8.58E-10       CGBO    = 1E-12
+CJ      = 9.465842E-4    PB      = 0.8            MJ      = 0.3722711
+CJSW    = 1.90832E-10    PBSW    = 0.8            MJSW    = 0.1366398
+CJSWG   = 3.3E-10        PBSWG   = 0.8            MJSWG   = 0.1366398
+CF      = 0              PVTH0   = -4.904276E-3   PRDSW   = -0.840458
+PK2     = 1.983844E-3    WKETA   = -1.794821E-3   LKETA   = -3.436309E-3
+PU0     = -3.6758958     PUA     = -4.70421E-11   PUB     = 8.241174E-24
+PVSAT   = 1.61878E3      PETA0   = 1E-4           PKETA   = -1.374594E-3    )
*
.MODEL PMOS PMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 4.1E-9
+XJ      = 1E-7           NCH     = 4.1589E17      VTH0    = -0.3901812
+K1      = 0.5723512      K2      = 0.024177       K3      = 0.1578539
+K3B     = 4.2732669      W0      = 1E-6           NLX     = 1.121486E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 0.6119889      DVT1    = 0.2499582      DVT2    = 0.1
+U0      = 112.2285112    UA      = 1.425392E-9    UB      = 1.16772E-21
+UC      = -1E-10         VSAT    = 1.087139E5     A0      = 1.5950482
+AGS     = 0.3203279      B0      = 4.957218E-7    B1      = 1.527303E-6
+KETA    = 0.0275656      A1      = 0.3799265      A2      = 0.432073
+RDSW    = 199.0599687    PRWG    = 0.5            PRWB    = -0.4953546
+WR      = 1              WINT    = 0              LINT    = 2.940415E-8
+         DWG     = -3.06329E-8
+DWB     = -7.685822E-9   VOFF    = -0.0937004     NFACTOR = 2
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 1.291671E-4    ETAB    = -2.161739E-4
+DSUB    = 3.645549E-4    PCLM    = 0.9284213      PDIBLC1 = 2.836414E-3
+PDIBLC2 = -8.750635E-6   PDIBLCB = -1E-3          DROUT   = 1.827199E-4
+PSCBE1  = 8E10           PSCBE2  = 8.26364E-10    PVAG    = 0.0202145
+DELTA   = 0.01           RSH     = 8.1            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 7.82E-10       CGSO    = 7.82E-10       CGBO    = 1E-12
+CJ      = 1.169586E-3    PB      = 0.8600389      MJ      = 0.4153558
+CJSW    = 2.172584E-10   PBSW    = 0.8            MJSW    = 0.3186705
+CJSWG   = 4.22E-10       PBSWG   = 0.8            MJSWG   = 0.3186705
+CF      = 0              PVTH0   = 1.231752E-3    PRDSW   = 9.5225138
+PK2     = 1.102104E-3    WKETA   = 0.0132876      LKETA   = -2.410443E-3
+PU0     = -1.5247633     PUA     = -5.27446E-11   PUB     = 1E-21
+PVSAT   = 50             PETA0   = 7.202744E-5    PKETA   = -1.607078E-3    )
*
